// Copyright (c) 2023 Beijing Institute of Open Source Chip
// common is licensed under Mulan PSL v2.
// You can use this software according to the terms and conditions of the Mulan PSL v2.
// You may obtain a copy of Mulan PSL v2 at:
//             http://license.coscl.org.cn/MulanPSL2
// THIS SOFTWARE IS PROVIDED ON AN "AS IS" BASIS, WITHOUT WARRANTIES OF ANY KIND,
// EITHER EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO NON-INFRINGEMENT,
// MERCHANTABILITY OR FIT FOR A PARTICULAR PURPOSE.
// See the Mulan PSL v2 for more details.

`ifndef INC_TEST_BASE_SV
`define INC_TEST_BASE_SV

class TestBase;
  string name;

  extern function new(string name = "test_base");
  extern task test_reset_register();
  extern task test_irq();
endclass

function TestBase::new(string name);
  this.name = name;
endfunction

task TestBase::test_reset_register();
  $display("=== [test reset register] ===");
endtask

task TestBase::test_irq();
  $display("=== [test irq] ===");
endtask

`endif
